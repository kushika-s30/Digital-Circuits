Half adder 
