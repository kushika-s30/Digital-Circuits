Half Adder 
